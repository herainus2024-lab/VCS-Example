`timescale 1ns/1ps

// ============================================================================
// UVM Top Testbench
// 顶层测试平台，实例化 DUT 并启动 UVM 测试
// ============================================================================
module tb_top;
  
  // 导入 UVM 和测试 package
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import multiplier_pkg::*;
  
  // ========================================================================
  // 时钟和复位
  // ========================================================================
  logic clk;
  logic rst_n;
  
  // 时钟生成 - 50MHz (周期 20ns)
  initial begin
    clk = 0;
    forever #10 clk = ~clk;
  end
  
  // 复位生成
  initial begin
    rst_n = 0;
    #50;
    rst_n = 1;
  end
  
  // ========================================================================
  // 接口实例化
  // ========================================================================
  multiplier_if aif(clk);
  
  // ========================================================================
  // DUT 实例化 (16-bit multiplier)
  // ========================================================================
  multiplier dut (
    .clk  (clk),
    .in1  (aif.in1),
    .in2  (aif.in2),
    .out  (aif.out)
  );
  
  // ========================================================================
  // 波形转储
  // ========================================================================
  initial begin
    // 支持 VCS/Verdi 波形
    `ifdef VCS
      $fsdbDumpfile("multiplier_uvm.fsdb");
      $fsdbDumpvars(0, tb_top);
      $fsdbDumpMDA();
    `endif
    
    // 支持其他仿真器
    `ifdef DUMP_VCD
      $dumpfile("multiplier_uvm.vcd");
      $dumpvars(0, tb_top);
    `endif
  end
  
  // ========================================================================
  // UVM 配置和启动
  // ========================================================================
  initial begin
    // 将接口传递给 UVM config_db
    uvm_config_db#(virtual multiplier_if)::set(null, "*", "vif", aif);
    
    // 设置超时时间
    uvm_top.set_timeout(10ms, 0);
    
    // 启动 UVM 测试
    run_test();
  end
  
  // ========================================================================
  // 仿真时间限制（安全措施）
  // ========================================================================
  initial begin
    #1000000;  // 1ms 超时
    `uvm_fatal("TIMEOUT", "Simulation timeout!")
  end

endmodule : tb_top
